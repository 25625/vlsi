`timescale 1ns / 1ns
module orgate(c,a,b);
input a,b;
output c;
or(c,a,b);
endmodule