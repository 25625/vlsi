`timescale 1ns / 1ns
module norgate(c,a,b);
input a,b;
output c;
and(c,a,b);
endmodule