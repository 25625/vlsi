`timescale 1ns / 1ps

module nandgate(c,a,b);
input a,b;
output c;
nand(c,a,b);
endmodule
