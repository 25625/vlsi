`timescale 1ns / 1ns
module andgate(c,a,b);
input a,b;
output c;
and(c,a,b);
endmodule`timescale 1ns / 1ns
